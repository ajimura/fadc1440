-- megafunction wizard: %ALTIOBUF%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altiobuf_out 

-- ============================================================
-- File Name: Obuf.vhd
-- Megafunction Name(s):
-- 			altiobuf_out
--
-- Simulation Library Files(s):
-- 			cycloneive
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 14.0.0 Build 200 06/17/2014 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus II License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


--altiobuf_out CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" ENABLE_BUS_HOLD="FALSE" LEFT_SHIFT_SERIES_TERMINATION_CONTROL="FALSE" NUMBER_OF_CHANNELS=2 OPEN_DRAIN_OUTPUT="FALSE" PSEUDO_DIFFERENTIAL_MODE="FALSE" USE_DIFFERENTIAL_MODE="FALSE" USE_OE="TRUE" USE_TERMINATION_CONTROL="FALSE" datain dataout oe
--VERSION_BEGIN 14.0 cbx_altiobuf_out 2014:06:17:18:06:03:SJ cbx_mgl 2014:06:17:18:10:38:SJ cbx_stratixiii 2014:06:17:18:06:03:SJ cbx_stratixv 2014:06:17:18:06:03:SJ  VERSION_END

 LIBRARY cycloneive;
 USE cycloneive.all;

--synthesis_resources = cycloneive_io_obuf 2 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  Obuf_iobuf_out_e5t IS 
	 PORT 
	 ( 
		 datain	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 dataout	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 oe	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0) := (OTHERS => '1')
	 ); 
 END Obuf_iobuf_out_e5t;

 ARCHITECTURE RTL OF Obuf_iobuf_out_e5t IS

	 SIGNAL  wire_obufa_i	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_obufa_o	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_obufa_oe	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  oe_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 COMPONENT  cycloneive_io_obuf
	 GENERIC 
	 (
		bus_hold	:	STRING := "false";
		open_drain_output	:	STRING := "false";
		lpm_type	:	STRING := "cycloneive_io_obuf"
	 );
	 PORT
	 ( 
		i	:	IN STD_LOGIC := '0';
		o	:	OUT STD_LOGIC;
		obar	:	OUT STD_LOGIC;
		oe	:	IN STD_LOGIC := '1';
		seriesterminationcontrol	:	IN STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	dataout <= wire_obufa_o;
	oe_w <= oe;
	wire_obufa_i <= datain;
	wire_obufa_oe <= oe_w;
	loop0 : FOR i IN 0 TO 1 GENERATE 
	  obufa :  cycloneive_io_obuf
	  GENERIC MAP (
		bus_hold => "false",
		open_drain_output => "false"
	  )
	  PORT MAP ( 
		i => wire_obufa_i(i),
		o => wire_obufa_o(i),
		oe => wire_obufa_oe(i)
	  );
	END GENERATE loop0;

 END RTL; --Obuf_iobuf_out_e5t
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Obuf IS
	PORT
	(
		datain		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		oe		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		dataout		: OUT STD_LOGIC_VECTOR (1 DOWNTO 0)
	);
END Obuf;


ARCHITECTURE RTL OF obuf IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (1 DOWNTO 0);



	COMPONENT Obuf_iobuf_out_e5t
	PORT (
			datain	: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
			oe	: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
			dataout	: OUT STD_LOGIC_VECTOR (1 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	dataout    <= sub_wire0(1 DOWNTO 0);

	Obuf_iobuf_out_e5t_component : Obuf_iobuf_out_e5t
	PORT MAP (
		datain => datain,
		oe => oe,
		dataout => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: enable_bus_hold STRING "FALSE"
-- Retrieval info: CONSTANT: left_shift_series_termination_control STRING "FALSE"
-- Retrieval info: CONSTANT: number_of_channels NUMERIC "2"
-- Retrieval info: CONSTANT: open_drain_output STRING "FALSE"
-- Retrieval info: CONSTANT: pseudo_differential_mode STRING "FALSE"
-- Retrieval info: CONSTANT: use_differential_mode STRING "FALSE"
-- Retrieval info: CONSTANT: use_oe STRING "TRUE"
-- Retrieval info: CONSTANT: use_termination_control STRING "FALSE"
-- Retrieval info: USED_PORT: datain 0 0 2 0 INPUT NODEFVAL "datain[1..0]"
-- Retrieval info: USED_PORT: dataout 0 0 2 0 OUTPUT NODEFVAL "dataout[1..0]"
-- Retrieval info: USED_PORT: oe 0 0 2 0 INPUT NODEFVAL "oe[1..0]"
-- Retrieval info: CONNECT: @datain 0 0 2 0 datain 0 0 2 0
-- Retrieval info: CONNECT: @oe 0 0 2 0 oe 0 0 2 0
-- Retrieval info: CONNECT: dataout 0 0 2 0 @dataout 0 0 2 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL Obuf.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Obuf.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Obuf.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Obuf.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Obuf_inst.vhd FALSE
-- Retrieval info: LIB_FILE: cycloneive
