    Mac OS X            	   2   �      �                                      ATTR       �   �                     �     !com.apple.genstore.origposixname ChBufManPeak.vhd